IXA00366430 00:25:b3:ca:5b:96 10.243.18.216 /BLANK/ROOT/PATH
IXA00342559 00:22:64:33:59:37 10.243.18.123 /BLANK/ROOT/PATH
IXA00342560 00:23:7D:1B:AE:A6 10.243.18.131 /BLANK/ROOT/PATH
IXA00342561 00:23:7D:1B:B1:DC 10.243.18.137 /BLANK/ROOT/PATH
IXA00366017 18:A9:05:EF:BC:53 10.243.18.192 /BLANK/ROOT/PATH
IXA00366508 00:09:6B:07:F0:FB 10.243.18.219 /BLANK/ROOT/PATH
IXA00372771 D0:67:E5:76:B9:77 10.243.18.244 /BLANK/ROOT/PATH
IXA00366014 00:13:20:F8:83:4B 10.243.18.189 /BLANK/ROOT/PATH
IXA00383418 00:13:20:FD:DF:3F 10.243.18.195 /BLANK/ROOT/PATH
IXA00371572 00:1e:67:2c:77:9f 10.243.18.108 /BLANK/ROOT/PATH
IXA00369888 00:E0:86:18:3A:A5 10.243.18.169 /BLANK/ROOT/PATH
IXA00369889 00:E0:86:17:00:32 10.243.18.221 /BLANK/ROOT/PATH
IXA00369890 00:e0:86:1b:bf:36 10.243.18.127 /BLANK/ROOT/PATH
IXA00369703 70:71:BC:DC:D0:1B 10.243.18.230 /BLANK/ROOT/PATH
IXA00369304 78:2B:CB:AF:1E:C1 10.243.18.199 /BLANK/ROOT/PATH
IXA00383377 00:13:20:FD:DF:08 10.243.18.139 /BLANK/ROOT/PATH
IXA00370123 00:E0:86:18:26:58 10.243.18.117 /BLANK/ROOT/PATH
IXA00370127 00:E0:86:18:21:4E 10.243.18.205 /BLANK/ROOT/PATH
IXA00370137 00:E0:86:16:C4:2E 10.243.18.51 /BLANK/ROOT/PATH
IXA00370141 00:E0:86:18:3A:9A 10.243.18.180 /BLANK/ROOT/PATH
IXA00381213 00:01:80:7D:F1:8F 10.243.18.81 /BLANK/ROOT/PATH
IXA00372626 00:30:48:B3:56:38 10.243.18.125 /BLANK/ROOT/PATH
IXA00382054 08:00:27:F3:F1:AB 10.243.18.162 /BLANK/ROOT/PATH
IXA00380890 00:11:22:23:24:25 10.243.18.97 /BLANK/ROOT/PATH
IXA00371002 38:60:77:12:50:c3 10.243.18.251 /BLANK/ROOT/PATH
IXA00380891 00:27:23:67:86:5b 10.243.18.156 /BLANK/ROOT/PATH
IXA00369786 00:80:a3:8c:81:6d 10.243.18.98 /BLANK/ROOT/PATH
IXA00383203 00:1e:67:56:b8:3a 10.243.18.154 /BLANK/ROOT/PATH
IXA00370130 00:E0:86:18:3A:9F 10.243.18.129 /BLANK/ROOT/PATH
IXA00382061 ec:a8:6b:f4:4e:aa 10.243.18.90 /BLANK/ROOT/PATH
IXA00372149 00:26:22:67:86:5B 10.243.18.133 /BLANK/ROOT/PATH
IXA00365684 00:15:17:be:28:5e 10.243.18.232 /BLANK/ROOT/PATH
IXA00366184 00:15:17:95:09:9d 10.243.18.181 /BLANK/ROOT/PATH
IXA00370133 00:E0:86:16:C4:36 10.243.18.248 /BLANK/ROOT/PATH
IXA00370385 00:E0:86:18:3B:78 10.243.18.159 /BLANK/ROOT/PATH
IXA00370839 E0:69:95:EB:75:CD 10.243.18.233 /BLANK/ROOT/PATH
IXA00379666 00:1E:67:43:4A:3A 10.243.18.106 /BLANK/ROOT/PATH
IXA00379966 68:05:CA:09:63:E8 10.243.18.66 /BLANK/ROOT/PATH
IXA00372507 00:15:17:BE:26:DB 10.243.18.110 /BLANK/ROOT/PATH
IXA00379576 E0:69:95:D3:0D:1B 10.243.18.103 /BLANK/ROOT/PATH
IXA00379771 00:e0:86:1b:bf:33 10.243.18.243 /BLANK/ROOT/PATH
IXA00370365 18:03:73:C6:EE:F1 10.243.18.165 /BLANK/ROOT/PATH
IXA00370367 18:03:73:C8:48:10 10.243.18.105 /BLANK/ROOT/PATH
IXA00382037 00:13:20:FD:D8:39 10.243.18.196 /BLANK/ROOT/PATH
IXA00382950 00:13:20:FD:DC:BA 10.243.18.253 /BLANK/ROOT/PATH
IXA00365421 00:15:17:DC:C6:5E 10.243.18.148 /BLANK/ROOT/PATH
IXA00372153 E0:69:95:D3:05:47 10.243.18.87 /BLANK/ROOT/PATH
IXA00383341 00:13:20:FD:DE:17 10.243.18.23 /BLANK/ROOT/PATH
IXA00372516 38:60:77:12:74:C0 10.243.18.254 /BLANK/ROOT/PATH
IXA00380742 68:05:ca:08:6b:e4 10.243.18.99 /BLANK/ROOT/PATH
IXA00378137 00:1e:67:3c:a3:7c 10.243.18.200 /BLANK/ROOT/PATH
IXA00380640 00:13:20:fd:09:48 10.243.18.150 /BLANK/ROOT/PATH
IXA00382137 00:13:20:FD:D8:E1 10.243.18.172 /BLANK/ROOT/PATH
IXA00370838 E0:69:95:E4:F6:D2 10.243.18.161 /BLANK/ROOT/PATH
IXA00383422 00:13:20:FD:DE:64 10.243.18.231 /BLANK/ROOT/PATH
IXA00380387 90:2B:34:5B:21:A8 10.243.18.223 /BLANK/ROOT/PATH
IXA00380551 90:2B:34:5B:1B:E6 10.243.18.14 /BLANK/ROOT/PATH
IXA00369959 38:60:77:12:87:AE 10.243.18.93 /BLANK/ROOT/PATH
IXA00380743 00:1B:21:00:6C:45 10.243.18.134 /BLANK/ROOT/PATH
IXA00365672 00:15:17:C5:1E:08 10.243.18.170 /BLANK/ROOT/PATH
IXA00381585 00:13:20:FD:D3:C6 10.243.18.166 /BLANK/ROOT/PATH
IXA00382138 00:13:20:FD:D8:1F 10.243.18.249 /BLANK/ROOT/PATH
IXA00368862 00:01:80:7C:9E:CD 10.243.18.53 /BLANK/ROOT/PATH
IXA00383755 00:13:20:FD:F3:80 10.243.18.115 /BLANK/ROOT/PATH
IXA00371944 38:60:77:12:8d:07 10.243.18.179 /BLANK/ROOT/PATH
IXA00372535 E0:69:95:EB:3D:06 10.243.18.118 /BLANK/ROOT/PATH
IXA00383081 00:13:20:FD:DC:B3 10.243.18.149 /BLANK/ROOT/PATH
IXA00372465 E0:69:95:EB:48:2E 10.243.18.140 /BLANK/ROOT/PATH
IXA00383732 00:13:20:FF:08:0E 10.243.18.160 /BLANK/ROOT/PATH
IXA00383754 00:13:20:FD:F3:5B 10.243.18.7 /BLANK/ROOT/PATH
IXA00383735 00:13:20:FD:F3:DA 10.243.18.143 /BLANK/ROOT/PATH
IXA00383021 00:13:20:fd:23:3d 10.243.18.5 /BLANK/ROOT/PATH
IXA00368470 00:15:17:a1:c2:7e 10.243.18.114 /BLANK/ROOT/PATH
IXA00378236 00:1B:21:4D:DF:D9 10.243.18.146 /BLANK/ROOT/PATH
